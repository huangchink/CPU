module shift(shift_type,shift_number,reg_data,shift_out);

input [1:0]shift_type;
input [4:0]shift_number;
input [31:0]reg_data;
output [31:0]shift_out;


reg [31:0]shift_out;
reg [31:0]temp;
reg [31:0]temp2,temp3;


always@(*)begin

temp=reg_data;
	case(shift_type)
		2'b00:
				shift_out=temp<<shift_number;
		2'b01:
				shift_out=temp>>shift_number;
		2'b10:begin
				case(shift_number)
				5'b00000:shift_out=reg_data;
				5'b00001:begin
							shift_out=temp>>1;
							shift_out[31]=reg_data[31];
							end
				5'b00010:begin
							shift_out=temp>>2;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							end
				5'b00011:begin
							shift_out=temp>>3;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							end
				5'b00100:begin
							shift_out=temp>>4;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							end
				5'b00101:begin
							shift_out=temp>>5;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							end
				5'b00110:begin
							shift_out=temp>>6;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							end
				5'b00111:begin
							shift_out=temp>>7;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							end
				5'b01000:begin
							shift_out=temp>>8;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							end
				5'b01001:begin
							shift_out=temp>>9;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							end
				5'b01010:begin
							shift_out=temp>>10;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							end
				5'b01011:begin
							shift_out=temp>>11;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							end
				5'b01100:begin
							shift_out=temp>>12;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							end
				5'b01101:begin
							shift_out=temp>>13;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							end
				5'b01110:begin
							shift_out=temp>>14;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							end
				5'b01111:begin
							shift_out=temp>>15;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							end
				5'b10000:begin
							shift_out=temp>>16;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							end
				5'b10001:begin
							shift_out=temp>>17;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							end
				5'b10010:begin
							shift_out=temp>>18;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							end
				5'b10011:begin
							shift_out=temp>>19;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							end
				5'b10100:begin
							shift_out=temp>>20;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							end
				5'b10101:begin
							shift_out=temp>>21;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							end
				5'b10110:begin
							shift_out=temp>>22;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							end
				5'b10111:begin
							shift_out=temp>>23;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							end
				5'b11000:begin
							shift_out=temp>>24;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							end
				5'b11001:begin
							shift_out=temp>>25;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							end
				5'b11010:begin
							shift_out=temp>>26;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							shift_out[6]=reg_data[31];
							end
				5'b11011:begin
							shift_out=temp>>27;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							shift_out[6]=reg_data[31];
							shift_out[5]=reg_data[31];
							end
				5'b11100:begin
							shift_out=temp>>28;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							shift_out[6]=reg_data[31];
							shift_out[5]=reg_data[31];
							shift_out[4]=reg_data[31];
							end
				5'b11101:begin
							shift_out=temp>>29;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							shift_out[6]=reg_data[31];
							shift_out[5]=reg_data[31];
							shift_out[4]=reg_data[31];
							shift_out[3]=reg_data[31];
							end		
				5'b11110:begin
							shift_out=temp>>30;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							shift_out[6]=reg_data[31];
							shift_out[5]=reg_data[31];
							shift_out[4]=reg_data[31];
							shift_out[3]=reg_data[31];
							shift_out[2]=reg_data[31];
							end	
				5'b11111:begin
							shift_out=temp>>31;
							shift_out[31]=reg_data[31];
							shift_out[30]=reg_data[31];
							shift_out[29]=reg_data[31];
							shift_out[28]=reg_data[31];
							shift_out[27]=reg_data[31];
							shift_out[26]=reg_data[31];
							shift_out[25]=reg_data[31];
							shift_out[24]=reg_data[31];
							shift_out[23]=reg_data[31];
							shift_out[22]=reg_data[31];
							shift_out[21]=reg_data[31];
							shift_out[20]=reg_data[31];
							shift_out[19]=reg_data[31];
							shift_out[18]=reg_data[31];
							shift_out[17]=reg_data[31];
							shift_out[16]=reg_data[31];
							shift_out[15]=reg_data[31];
							shift_out[14]=reg_data[31];
							shift_out[13]=reg_data[31];
							shift_out[12]=reg_data[31];
							shift_out[11]=reg_data[31];
							shift_out[10]=reg_data[31];
							shift_out[9]=reg_data[31];
							shift_out[8]=reg_data[31];
							shift_out[7]=reg_data[31];
							shift_out[6]=reg_data[31];
							shift_out[5]=reg_data[31];
							shift_out[4]=reg_data[31];
							shift_out[3]=reg_data[31];
							shift_out[2]=reg_data[31];
							end									
					endcase
				end
				
		2'b11:begin
				case(shift_type)
				5'b00000:shift_out=reg_data;
				5'b00001:begin
							shift_out=temp>>1;
							shift_out[31]=reg_data[0];
							end
				5'b00010:begin
							shift_out=temp>>2;
							shift_out[31]=reg_data[1];
							shift_out[30]=reg_data[0];
							end
				5'b00011:begin
							shift_out=temp>>3;
							shift_out[31]=reg_data[2];
							shift_out[30]=reg_data[1];
							shift_out[29]=reg_data[0];
							end
				5'b00100:begin
							shift_out=temp>>4;
							shift_out[31]=reg_data[3];
							shift_out[30]=reg_data[2];
							shift_out[29]=reg_data[1];
							shift_out[28]=reg_data[0];
							end
				5'b00101:begin
							shift_out=temp>>5;
							shift_out[31]=reg_data[4];
							shift_out[30]=reg_data[3];
							shift_out[29]=reg_data[2];
							shift_out[28]=reg_data[1];
							shift_out[27]=reg_data[0];
							end
				5'b00110:begin
							shift_out=temp>>6;
							shift_out[31]=reg_data[5];
							shift_out[30]=reg_data[4];
							shift_out[29]=reg_data[3];
							shift_out[28]=reg_data[2];
							shift_out[27]=reg_data[1];
							shift_out[26]=reg_data[0];
							end
				5'b00111:begin
							shift_out=temp>>7;
							shift_out[31]=reg_data[6];
							shift_out[30]=reg_data[5];
							shift_out[29]=reg_data[4];
							shift_out[28]=reg_data[3];
							shift_out[27]=reg_data[2];
							shift_out[26]=reg_data[1];
							shift_out[25]=reg_data[0];
							end
				5'b01000:begin
							shift_out=temp>>8;
							shift_out[31]=reg_data[7];
							shift_out[30]=reg_data[6];
							shift_out[29]=reg_data[5];
							shift_out[28]=reg_data[4];
							shift_out[27]=reg_data[3];
							shift_out[26]=reg_data[2];
							shift_out[25]=reg_data[1];
							shift_out[24]=reg_data[0];
							end
				5'b01001:begin
							shift_out=temp>>9;
							shift_out[31]=reg_data[8];
							shift_out[30]=reg_data[7];
							shift_out[29]=reg_data[6];
							shift_out[28]=reg_data[5];
							shift_out[27]=reg_data[4];
							shift_out[26]=reg_data[3];
							shift_out[25]=reg_data[2];
							shift_out[24]=reg_data[1];
							shift_out[23]=reg_data[0];
							end
				5'b01010:begin
							shift_out=temp>>10;
							shift_out[31]=reg_data[9];
							shift_out[30]=reg_data[8];
							shift_out[29]=reg_data[7];
							shift_out[28]=reg_data[6];
							shift_out[27]=reg_data[5];
							shift_out[26]=reg_data[4];
							shift_out[25]=reg_data[3];
							shift_out[24]=reg_data[2];
							shift_out[23]=reg_data[1];
							shift_out[22]=reg_data[0];
							end
				5'b01011:begin
							shift_out=temp>>11;
							shift_out[31]=reg_data[10];
							shift_out[30]=reg_data[9];
							shift_out[29]=reg_data[8];
							shift_out[28]=reg_data[7];
							shift_out[27]=reg_data[6];
							shift_out[26]=reg_data[5];
							shift_out[25]=reg_data[4];
							shift_out[24]=reg_data[3];
							shift_out[23]=reg_data[2];
							shift_out[22]=reg_data[1];
							shift_out[21]=reg_data[0];
							end
				5'b01100:begin
							shift_out=temp>>12;
							shift_out[31]=reg_data[11];
							shift_out[30]=reg_data[10];
							shift_out[29]=reg_data[9];
							shift_out[28]=reg_data[8];
							shift_out[27]=reg_data[7];
							shift_out[26]=reg_data[6];
							shift_out[25]=reg_data[5];
							shift_out[24]=reg_data[4];
							shift_out[23]=reg_data[3];
							shift_out[22]=reg_data[2];
							shift_out[21]=reg_data[1];
							shift_out[20]=reg_data[0];
							end
				5'b01101:begin
							shift_out=temp>>13;
							shift_out[31]=reg_data[12];
							shift_out[30]=reg_data[11];
							shift_out[29]=reg_data[10];
							shift_out[28]=reg_data[9];
							shift_out[27]=reg_data[8];
							shift_out[26]=reg_data[7];
							shift_out[25]=reg_data[6];
							shift_out[24]=reg_data[5];
							shift_out[23]=reg_data[4];
							shift_out[22]=reg_data[3];
							shift_out[21]=reg_data[2];
							shift_out[20]=reg_data[1];
							shift_out[19]=reg_data[0];
							end
				5'b01110:begin
							shift_out=temp>>14;
							shift_out[31]=reg_data[13];
							shift_out[30]=reg_data[12];
							shift_out[29]=reg_data[11];
							shift_out[28]=reg_data[10];
							shift_out[27]=reg_data[9];
							shift_out[26]=reg_data[8];
							shift_out[25]=reg_data[7];
							shift_out[24]=reg_data[6];
							shift_out[23]=reg_data[5];
							shift_out[22]=reg_data[4];
							shift_out[21]=reg_data[3];
							shift_out[20]=reg_data[2];
							shift_out[19]=reg_data[1];
							shift_out[18]=reg_data[0];
							end
				5'b01111:begin
							shift_out=temp>>15;
							shift_out[31]=reg_data[14];
							shift_out[30]=reg_data[13];
							shift_out[29]=reg_data[12];
							shift_out[28]=reg_data[11];
							shift_out[27]=reg_data[10];
							shift_out[26]=reg_data[9];
							shift_out[25]=reg_data[8];
							shift_out[24]=reg_data[7];
							shift_out[23]=reg_data[6];
							shift_out[22]=reg_data[5];
							shift_out[21]=reg_data[4];
							shift_out[20]=reg_data[3];
							shift_out[19]=reg_data[2];
							shift_out[18]=reg_data[1];
							shift_out[17]=reg_data[0];
							end
				5'b10000:begin
							shift_out=temp>>16;
							shift_out[31]=reg_data[15];
							shift_out[30]=reg_data[14];
							shift_out[29]=reg_data[13];
							shift_out[28]=reg_data[12];
							shift_out[27]=reg_data[11];
							shift_out[26]=reg_data[10];
							shift_out[25]=reg_data[9];
							shift_out[24]=reg_data[8];
							shift_out[23]=reg_data[7];
							shift_out[22]=reg_data[6];
							shift_out[21]=reg_data[5];
							shift_out[20]=reg_data[4];
							shift_out[19]=reg_data[3];
							shift_out[18]=reg_data[2];
							shift_out[17]=reg_data[1];
							shift_out[16]=reg_data[0];
							end
				5'b10001:begin
							shift_out=temp>>17;
							shift_out[31]=reg_data[16];
							shift_out[30]=reg_data[15];
							shift_out[29]=reg_data[14];
							shift_out[28]=reg_data[13];
							shift_out[27]=reg_data[12];
							shift_out[26]=reg_data[11];
							shift_out[25]=reg_data[10];
							shift_out[24]=reg_data[9];
							shift_out[23]=reg_data[8];
							shift_out[22]=reg_data[7];
							shift_out[21]=reg_data[6];
							shift_out[20]=reg_data[5];
							shift_out[19]=reg_data[4];
							shift_out[18]=reg_data[3];
							shift_out[17]=reg_data[2];
							shift_out[16]=reg_data[1];
							shift_out[15]=reg_data[0];
							end
				5'b10010:begin
							shift_out=temp>>18;
							shift_out[31]=reg_data[17];
							shift_out[30]=reg_data[16];
							shift_out[29]=reg_data[15];
							shift_out[28]=reg_data[14];
							shift_out[27]=reg_data[13];
							shift_out[26]=reg_data[12];
							shift_out[25]=reg_data[11];
							shift_out[24]=reg_data[10];
							shift_out[23]=reg_data[9];
							shift_out[22]=reg_data[8];
							shift_out[21]=reg_data[7];
							shift_out[20]=reg_data[6];
							shift_out[19]=reg_data[5];
							shift_out[18]=reg_data[4];
							shift_out[17]=reg_data[3];
							shift_out[16]=reg_data[2];
							shift_out[15]=reg_data[1];
							shift_out[14]=reg_data[0];
							end
				5'b10011:begin
							shift_out=temp>>19;
							shift_out[31]=reg_data[18];
							shift_out[30]=reg_data[17];
							shift_out[29]=reg_data[16];
							shift_out[28]=reg_data[15];
							shift_out[27]=reg_data[14];
							shift_out[26]=reg_data[13];
							shift_out[25]=reg_data[12];
							shift_out[24]=reg_data[11];
							shift_out[23]=reg_data[10];
							shift_out[22]=reg_data[9];
							shift_out[21]=reg_data[8];
							shift_out[20]=reg_data[7];
							shift_out[19]=reg_data[6];
							shift_out[18]=reg_data[5];
							shift_out[17]=reg_data[4];
							shift_out[16]=reg_data[3];
							shift_out[15]=reg_data[2];
							shift_out[14]=reg_data[1];
							shift_out[13]=reg_data[0];
							end
				5'b10100:begin
							shift_out=temp>>20;
							shift_out[31]=reg_data[19];
							shift_out[30]=reg_data[18];
							shift_out[29]=reg_data[17];
							shift_out[28]=reg_data[16];
							shift_out[27]=reg_data[15];
							shift_out[26]=reg_data[14];
							shift_out[25]=reg_data[13];
							shift_out[24]=reg_data[12];
							shift_out[23]=reg_data[11];
							shift_out[22]=reg_data[10];
							shift_out[21]=reg_data[9];
							shift_out[20]=reg_data[8];
							shift_out[19]=reg_data[7];
							shift_out[18]=reg_data[6];
							shift_out[17]=reg_data[5];
							shift_out[16]=reg_data[4];
							shift_out[15]=reg_data[3];
							shift_out[14]=reg_data[2];
							shift_out[13]=reg_data[1];
							shift_out[12]=reg_data[0];
							end
				5'b10101:begin
							shift_out=temp>>21;
							shift_out[31]=reg_data[20];
							shift_out[30]=reg_data[19];
							shift_out[29]=reg_data[18];
							shift_out[28]=reg_data[17];
							shift_out[27]=reg_data[16];
							shift_out[26]=reg_data[15];
							shift_out[25]=reg_data[14];
							shift_out[24]=reg_data[13];
							shift_out[23]=reg_data[12];
							shift_out[22]=reg_data[11];
							shift_out[21]=reg_data[10];
							shift_out[20]=reg_data[9];
							shift_out[19]=reg_data[8];
							shift_out[18]=reg_data[7];
							shift_out[17]=reg_data[6];
							shift_out[16]=reg_data[5];
							shift_out[15]=reg_data[4];
							shift_out[14]=reg_data[3];
							shift_out[13]=reg_data[2];
							shift_out[12]=reg_data[1];
							shift_out[11]=reg_data[0];
							end
				5'b10110:begin
							shift_out=temp>>22;
							shift_out[31]=reg_data[21];
							shift_out[30]=reg_data[20];
							shift_out[29]=reg_data[19];
							shift_out[28]=reg_data[18];
							shift_out[27]=reg_data[17];
							shift_out[26]=reg_data[16];
							shift_out[25]=reg_data[15];
							shift_out[24]=reg_data[14];
							shift_out[23]=reg_data[13];
							shift_out[22]=reg_data[12];
							shift_out[21]=reg_data[11];
							shift_out[20]=reg_data[10];
							shift_out[19]=reg_data[9];
							shift_out[18]=reg_data[8];
							shift_out[17]=reg_data[7];
							shift_out[16]=reg_data[6];
							shift_out[15]=reg_data[5];
							shift_out[14]=reg_data[4];
							shift_out[13]=reg_data[3];
							shift_out[12]=reg_data[2];
							shift_out[11]=reg_data[1];
							shift_out[10]=reg_data[0];
							end
				5'b10111:begin
							shift_out=temp>>23;
							shift_out[31]=reg_data[22];
							shift_out[30]=reg_data[21];
							shift_out[29]=reg_data[20];
							shift_out[28]=reg_data[19];
							shift_out[27]=reg_data[18];
							shift_out[26]=reg_data[17];
							shift_out[25]=reg_data[16];
							shift_out[24]=reg_data[15];
							shift_out[23]=reg_data[14];
							shift_out[22]=reg_data[13];
							shift_out[21]=reg_data[12];
							shift_out[20]=reg_data[11];
							shift_out[19]=reg_data[10];
							shift_out[18]=reg_data[9];
							shift_out[17]=reg_data[8];
							shift_out[16]=reg_data[7];
							shift_out[15]=reg_data[6];
							shift_out[14]=reg_data[5];
							shift_out[13]=reg_data[4];
							shift_out[12]=reg_data[3];
							shift_out[11]=reg_data[2];
							shift_out[10]=reg_data[1];
							shift_out[9]=reg_data[0];
							end
				5'b11000:begin
							shift_out=temp>>24;
							shift_out[31]=reg_data[23];
							shift_out[30]=reg_data[22];
							shift_out[29]=reg_data[21];
							shift_out[28]=reg_data[20];
							shift_out[27]=reg_data[19];
							shift_out[26]=reg_data[18];
							shift_out[25]=reg_data[17];
							shift_out[24]=reg_data[16];
							shift_out[23]=reg_data[15];
							shift_out[22]=reg_data[14];
							shift_out[21]=reg_data[13];
							shift_out[20]=reg_data[12];
							shift_out[19]=reg_data[11];
							shift_out[18]=reg_data[10];
							shift_out[17]=reg_data[9];
							shift_out[16]=reg_data[8];
							shift_out[15]=reg_data[7];
							shift_out[14]=reg_data[6];
							shift_out[13]=reg_data[5];
							shift_out[12]=reg_data[4];
							shift_out[11]=reg_data[3];
							shift_out[10]=reg_data[2];
							shift_out[9]=reg_data[1];
							shift_out[8]=reg_data[0];
							end
				5'b11001:begin
							shift_out=temp>>25;
							shift_out[31]=reg_data[24];
							shift_out[30]=reg_data[23];
							shift_out[29]=reg_data[22];
							shift_out[28]=reg_data[21];
							shift_out[27]=reg_data[20];
							shift_out[26]=reg_data[19];
							shift_out[25]=reg_data[18];
							shift_out[24]=reg_data[17];
							shift_out[23]=reg_data[16];
							shift_out[22]=reg_data[15];
							shift_out[21]=reg_data[14];
							shift_out[20]=reg_data[13];
							shift_out[19]=reg_data[12];
							shift_out[18]=reg_data[11];
							shift_out[17]=reg_data[10];
							shift_out[16]=reg_data[9];
							shift_out[15]=reg_data[8];
							shift_out[14]=reg_data[7];
							shift_out[13]=reg_data[6];
							shift_out[12]=reg_data[5];
							shift_out[11]=reg_data[4];
							shift_out[10]=reg_data[3];
							shift_out[9]=reg_data[2];
							shift_out[8]=reg_data[1];
							shift_out[7]=reg_data[0];
							end
				5'b11010:begin
							shift_out=temp>>26;
							shift_out[31]=reg_data[25];
							shift_out[30]=reg_data[24];
							shift_out[29]=reg_data[23];
							shift_out[28]=reg_data[22];
							shift_out[27]=reg_data[21];
							shift_out[26]=reg_data[20];
							shift_out[25]=reg_data[19];
							shift_out[24]=reg_data[18];
							shift_out[23]=reg_data[17];
							shift_out[22]=reg_data[16];
							shift_out[21]=reg_data[15];
							shift_out[20]=reg_data[14];
							shift_out[19]=reg_data[13];
							shift_out[18]=reg_data[12];
							shift_out[17]=reg_data[11];
							shift_out[16]=reg_data[10];
							shift_out[15]=reg_data[9];
							shift_out[14]=reg_data[8];
							shift_out[13]=reg_data[7];
							shift_out[12]=reg_data[6];
							shift_out[11]=reg_data[5];
							shift_out[10]=reg_data[4];
							shift_out[9]=reg_data[3];
							shift_out[8]=reg_data[2];
							shift_out[7]=reg_data[1];
							shift_out[6]=reg_data[0];
							end
				5'b11011:begin
							shift_out=temp>>27;
							shift_out[31]=reg_data[26];
							shift_out[30]=reg_data[25];
							shift_out[29]=reg_data[24];
							shift_out[28]=reg_data[23];
							shift_out[27]=reg_data[22];
							shift_out[26]=reg_data[21];
							shift_out[25]=reg_data[20];
							shift_out[24]=reg_data[19];
							shift_out[23]=reg_data[18];
							shift_out[22]=reg_data[17];
							shift_out[21]=reg_data[16];
							shift_out[20]=reg_data[15];
							shift_out[19]=reg_data[14];
							shift_out[18]=reg_data[13];
							shift_out[17]=reg_data[12];
							shift_out[16]=reg_data[11];
							shift_out[15]=reg_data[10];
							shift_out[14]=reg_data[9];
							shift_out[13]=reg_data[8];
							shift_out[12]=reg_data[7];
							shift_out[11]=reg_data[6];
							shift_out[10]=reg_data[5];
							shift_out[9]=reg_data[4];
							shift_out[8]=reg_data[3];
							shift_out[7]=reg_data[2];
							shift_out[6]=reg_data[1];
							shift_out[5]=reg_data[0];
							end
				5'b11100:begin
							shift_out=temp>>28;
							shift_out[31]=reg_data[27];
							shift_out[30]=reg_data[26];
							shift_out[29]=reg_data[25];
							shift_out[28]=reg_data[24];
							shift_out[27]=reg_data[23];
							shift_out[26]=reg_data[22];
							shift_out[25]=reg_data[21];
							shift_out[24]=reg_data[20];
							shift_out[23]=reg_data[19];
							shift_out[22]=reg_data[18];
							shift_out[21]=reg_data[17];
							shift_out[20]=reg_data[16];
							shift_out[19]=reg_data[15];
							shift_out[18]=reg_data[14];
							shift_out[17]=reg_data[13];
							shift_out[16]=reg_data[12];
							shift_out[15]=reg_data[11];
							shift_out[14]=reg_data[10];
							shift_out[13]=reg_data[9];
							shift_out[12]=reg_data[8];
							shift_out[11]=reg_data[7];
							shift_out[10]=reg_data[6];
							shift_out[9]=reg_data[5];
							shift_out[8]=reg_data[4];
							shift_out[7]=reg_data[3];
							shift_out[6]=reg_data[2];
							shift_out[5]=reg_data[1];
							shift_out[4]=reg_data[0];
							end
				5'b11101:begin
							shift_out=temp>>29;
							shift_out[31]=reg_data[28];
							shift_out[30]=reg_data[27];
							shift_out[29]=reg_data[26];
							shift_out[28]=reg_data[25];
							shift_out[27]=reg_data[24];
							shift_out[26]=reg_data[23];
							shift_out[25]=reg_data[22];
							shift_out[24]=reg_data[21];
							shift_out[23]=reg_data[20];
							shift_out[22]=reg_data[19];
							shift_out[21]=reg_data[18];
							shift_out[20]=reg_data[17];
							shift_out[19]=reg_data[16];
							shift_out[18]=reg_data[15];
							shift_out[17]=reg_data[14];
							shift_out[16]=reg_data[13];
							shift_out[15]=reg_data[12];
							shift_out[14]=reg_data[11];
							shift_out[13]=reg_data[10];
							shift_out[12]=reg_data[9];
							shift_out[11]=reg_data[8];
							shift_out[10]=reg_data[7];
							shift_out[9]=reg_data[6];
							shift_out[8]=reg_data[5];
							shift_out[7]=reg_data[4];
							shift_out[6]=reg_data[3];
							shift_out[5]=reg_data[2];
							shift_out[4]=reg_data[1];
							shift_out[3]=reg_data[0];
							end		
				5'b11110:begin
							shift_out=temp>>30;
							shift_out[31]=reg_data[29];
							shift_out[30]=reg_data[28];
							shift_out[29]=reg_data[27];
							shift_out[28]=reg_data[26];
							shift_out[27]=reg_data[25];
							shift_out[26]=reg_data[24];
							shift_out[25]=reg_data[23];
							shift_out[24]=reg_data[22];
							shift_out[23]=reg_data[21];
							shift_out[22]=reg_data[20];
							shift_out[21]=reg_data[19];
							shift_out[20]=reg_data[18];
							shift_out[19]=reg_data[17];
							shift_out[18]=reg_data[16];
							shift_out[17]=reg_data[15];
							shift_out[16]=reg_data[14];
							shift_out[15]=reg_data[13];
							shift_out[14]=reg_data[12];
							shift_out[13]=reg_data[11];
							shift_out[12]=reg_data[10];
							shift_out[11]=reg_data[9];
							shift_out[10]=reg_data[8];
							shift_out[9]=reg_data[7];
							shift_out[8]=reg_data[6];
							shift_out[7]=reg_data[5];
							shift_out[6]=reg_data[4];
							shift_out[5]=reg_data[3];
							shift_out[4]=reg_data[2];
							shift_out[3]=reg_data[1];
							shift_out[2]=reg_data[0];
							end	
				5'b11111:begin
							shift_out=temp>>31;
							shift_out[31]=reg_data[30];
							shift_out[30]=reg_data[29];
							shift_out[29]=reg_data[28];
							shift_out[28]=reg_data[27];
							shift_out[27]=reg_data[26];
							shift_out[26]=reg_data[25];
							shift_out[25]=reg_data[24];
							shift_out[24]=reg_data[23];
							shift_out[23]=reg_data[22];
							shift_out[22]=reg_data[21];
							shift_out[21]=reg_data[20];
							shift_out[20]=reg_data[19];
							shift_out[19]=reg_data[18];
							shift_out[18]=reg_data[17];
							shift_out[17]=reg_data[16];
							shift_out[16]=reg_data[15];
							shift_out[15]=reg_data[14];
							shift_out[14]=reg_data[13];
							shift_out[13]=reg_data[12];
							shift_out[12]=reg_data[11];
							shift_out[11]=reg_data[10];
							shift_out[10]=reg_data[9];
							shift_out[9]=reg_data[8];
							shift_out[8]=reg_data[7];
							shift_out[7]=reg_data[6];
							shift_out[6]=reg_data[5];
							shift_out[5]=reg_data[4];
							shift_out[4]=reg_data[3];
							shift_out[3]=reg_data[2];
							shift_out[2]=reg_data[1];	
							shift_out[1]=reg_data[0];	
							end									
					endcase
				end
		 
	endcase
end
endmodule





 
 


