module rotate(immediate_in,rotate_immediate_out);

input [11:0]immediate_in;
output reg[31:0]rotate_immediate_out;

reg 	[31:0]extend_immediate_in;
reg 	[31:0]temp;


always@(*)begin

temp=32'b0;
extend_immediate_in=temp+immediate_in[7:0];
temp=extend_immediate_in;
	case(immediate_in[11:8])
	4'b0000:rotate_immediate_out=extend_immediate_in;
	4'b0001:begin
			  rotate_immediate_out=temp>>2;
			  rotate_immediate_out[31]=extend_immediate_in[1];
			  rotate_immediate_out[30]=extend_immediate_in[0];
			  end
	4'b0010:begin
			  rotate_immediate_out=temp>>4;
			  rotate_immediate_out[31]=extend_immediate_in[3];
			  rotate_immediate_out[30]=extend_immediate_in[2];
			  rotate_immediate_out[29]=extend_immediate_in[1];
			  rotate_immediate_out[28]=extend_immediate_in[0];
			  end
	4'b0011:begin
			  rotate_immediate_out=temp>>6;
			  rotate_immediate_out[31]=extend_immediate_in[5];
			  rotate_immediate_out[30]=extend_immediate_in[4];
			  rotate_immediate_out[29]=extend_immediate_in[3];
			  rotate_immediate_out[28]=extend_immediate_in[2];
			  rotate_immediate_out[27]=extend_immediate_in[1];
			  rotate_immediate_out[26]=extend_immediate_in[0];
			  end
	4'b0100:begin
			  rotate_immediate_out=temp>>8;
			  rotate_immediate_out[31]=extend_immediate_in[7];
			  rotate_immediate_out[30]=extend_immediate_in[6];
			  rotate_immediate_out[29]=extend_immediate_in[5];
			  rotate_immediate_out[28]=extend_immediate_in[4];
			  rotate_immediate_out[27]=extend_immediate_in[3];
			  rotate_immediate_out[26]=extend_immediate_in[2];
			  rotate_immediate_out[25]=extend_immediate_in[1];
			  rotate_immediate_out[24]=extend_immediate_in[0];
			  end
	4'b0101:begin
			  rotate_immediate_out=temp>>10;
			  rotate_immediate_out[31]=extend_immediate_in[9];
			  rotate_immediate_out[30]=extend_immediate_in[8];
			  rotate_immediate_out[29]=extend_immediate_in[7];
			  rotate_immediate_out[28]=extend_immediate_in[6];
			  rotate_immediate_out[27]=extend_immediate_in[5];
			  rotate_immediate_out[26]=extend_immediate_in[4];
			  rotate_immediate_out[25]=extend_immediate_in[3];
			  rotate_immediate_out[24]=extend_immediate_in[2];
			  rotate_immediate_out[23]=extend_immediate_in[1];
			  rotate_immediate_out[22]=extend_immediate_in[0];
			  end
	4'b0110:begin
			  rotate_immediate_out=temp>>12;
			  rotate_immediate_out[31]=extend_immediate_in[11];
			  rotate_immediate_out[30]=extend_immediate_in[10];
			  rotate_immediate_out[29]=extend_immediate_in[9];
			  rotate_immediate_out[28]=extend_immediate_in[8];
			  rotate_immediate_out[27]=extend_immediate_in[7];
			  rotate_immediate_out[26]=extend_immediate_in[6];
			  rotate_immediate_out[25]=extend_immediate_in[5];
			  rotate_immediate_out[24]=extend_immediate_in[4];
			  rotate_immediate_out[23]=extend_immediate_in[3];
			  rotate_immediate_out[22]=extend_immediate_in[2];
			  rotate_immediate_out[21]=extend_immediate_in[1];
			  rotate_immediate_out[20]=extend_immediate_in[0];
			  end
	4'b0111:begin
			  rotate_immediate_out=temp>>14;
			  rotate_immediate_out[31]=extend_immediate_in[13];
			  rotate_immediate_out[30]=extend_immediate_in[12];
			  rotate_immediate_out[29]=extend_immediate_in[11];
			  rotate_immediate_out[28]=extend_immediate_in[10];
			  rotate_immediate_out[27]=extend_immediate_in[9];
			  rotate_immediate_out[26]=extend_immediate_in[8];
			  rotate_immediate_out[25]=extend_immediate_in[7];
			  rotate_immediate_out[24]=extend_immediate_in[6];
			  rotate_immediate_out[23]=extend_immediate_in[5];
			  rotate_immediate_out[22]=extend_immediate_in[4];
			  rotate_immediate_out[21]=extend_immediate_in[3];
			  rotate_immediate_out[20]=extend_immediate_in[2];
			  rotate_immediate_out[19]=extend_immediate_in[1];
			  rotate_immediate_out[18]=extend_immediate_in[0];
			  end
	4'b1000:begin
			  rotate_immediate_out=temp>>16;
			  rotate_immediate_out[31]=extend_immediate_in[15];
			  rotate_immediate_out[30]=extend_immediate_in[14];
			  rotate_immediate_out[29]=extend_immediate_in[13];
			  rotate_immediate_out[28]=extend_immediate_in[12];
			  rotate_immediate_out[27]=extend_immediate_in[11];
			  rotate_immediate_out[26]=extend_immediate_in[10];
			  rotate_immediate_out[25]=extend_immediate_in[9];
			  rotate_immediate_out[24]=extend_immediate_in[8];
			  rotate_immediate_out[23]=extend_immediate_in[7];
			  rotate_immediate_out[22]=extend_immediate_in[6];
			  rotate_immediate_out[21]=extend_immediate_in[5];
			  rotate_immediate_out[20]=extend_immediate_in[4];
			  rotate_immediate_out[19]=extend_immediate_in[3];
			  rotate_immediate_out[18]=extend_immediate_in[2];
			  rotate_immediate_out[17]=extend_immediate_in[1];
			  rotate_immediate_out[16]=extend_immediate_in[0];
			  end
	4'b1001:begin
			  rotate_immediate_out=temp>>18;
			  rotate_immediate_out[31]=extend_immediate_in[17];
			  rotate_immediate_out[30]=extend_immediate_in[16];
			  rotate_immediate_out[29]=extend_immediate_in[15];
			  rotate_immediate_out[28]=extend_immediate_in[14];
			  rotate_immediate_out[27]=extend_immediate_in[13];
			  rotate_immediate_out[26]=extend_immediate_in[12];
			  rotate_immediate_out[25]=extend_immediate_in[11];
			  rotate_immediate_out[24]=extend_immediate_in[10];
			  rotate_immediate_out[23]=extend_immediate_in[9];
			  rotate_immediate_out[22]=extend_immediate_in[8];
			  rotate_immediate_out[21]=extend_immediate_in[7];
			  rotate_immediate_out[20]=extend_immediate_in[6];
			  rotate_immediate_out[19]=extend_immediate_in[5];
			  rotate_immediate_out[18]=extend_immediate_in[4];
			  rotate_immediate_out[17]=extend_immediate_in[3];
			  rotate_immediate_out[16]=extend_immediate_in[2];
			  rotate_immediate_out[15]=extend_immediate_in[1];
			  rotate_immediate_out[14]=extend_immediate_in[0];
			  end
	4'b1010:begin
			  rotate_immediate_out=temp>>20;
			  rotate_immediate_out[31]=extend_immediate_in[19];
			  rotate_immediate_out[30]=extend_immediate_in[18];
			  rotate_immediate_out[29]=extend_immediate_in[17];
			  rotate_immediate_out[28]=extend_immediate_in[16];
			  rotate_immediate_out[27]=extend_immediate_in[15];
			  rotate_immediate_out[26]=extend_immediate_in[14];
			  rotate_immediate_out[25]=extend_immediate_in[13];
			  rotate_immediate_out[24]=extend_immediate_in[12];
			  rotate_immediate_out[23]=extend_immediate_in[11];
			  rotate_immediate_out[22]=extend_immediate_in[10];
			  rotate_immediate_out[21]=extend_immediate_in[9];
			  rotate_immediate_out[20]=extend_immediate_in[8];
			  rotate_immediate_out[19]=extend_immediate_in[7];
			  rotate_immediate_out[18]=extend_immediate_in[6];
			  rotate_immediate_out[17]=extend_immediate_in[5];
			  rotate_immediate_out[16]=extend_immediate_in[4];
			  rotate_immediate_out[15]=extend_immediate_in[3];
			  rotate_immediate_out[14]=extend_immediate_in[2];
			  rotate_immediate_out[13]=extend_immediate_in[1];
			  rotate_immediate_out[12]=extend_immediate_in[0];
			  end
	4'b1011:begin
			  rotate_immediate_out=temp>>22;
			  rotate_immediate_out[31]=extend_immediate_in[21];
			  rotate_immediate_out[30]=extend_immediate_in[20];
			  rotate_immediate_out[29]=extend_immediate_in[19];
			  rotate_immediate_out[28]=extend_immediate_in[18];
			  rotate_immediate_out[27]=extend_immediate_in[17];
			  rotate_immediate_out[26]=extend_immediate_in[16];
			  rotate_immediate_out[25]=extend_immediate_in[15];
			  rotate_immediate_out[24]=extend_immediate_in[14];
			  rotate_immediate_out[23]=extend_immediate_in[13];
			  rotate_immediate_out[22]=extend_immediate_in[12];
			  rotate_immediate_out[21]=extend_immediate_in[11];
			  rotate_immediate_out[20]=extend_immediate_in[10];
			  rotate_immediate_out[19]=extend_immediate_in[9];
			  rotate_immediate_out[18]=extend_immediate_in[8];
			  rotate_immediate_out[17]=extend_immediate_in[7];
			  rotate_immediate_out[16]=extend_immediate_in[6];
			  rotate_immediate_out[15]=extend_immediate_in[5];
			  rotate_immediate_out[14]=extend_immediate_in[4];
			  rotate_immediate_out[13]=extend_immediate_in[3];
			  rotate_immediate_out[12]=extend_immediate_in[2];
			  rotate_immediate_out[11]=extend_immediate_in[1];
			  rotate_immediate_out[10]=extend_immediate_in[0];
			  end
	4'b1100:begin
			  rotate_immediate_out=temp>>24;
			  rotate_immediate_out[31]=extend_immediate_in[23];
			  rotate_immediate_out[30]=extend_immediate_in[22];
			  rotate_immediate_out[29]=extend_immediate_in[21];
			  rotate_immediate_out[28]=extend_immediate_in[20];
			  rotate_immediate_out[27]=extend_immediate_in[19];
			  rotate_immediate_out[26]=extend_immediate_in[18];
			  rotate_immediate_out[25]=extend_immediate_in[17];
			  rotate_immediate_out[24]=extend_immediate_in[16];
			  rotate_immediate_out[23]=extend_immediate_in[15];
			  rotate_immediate_out[22]=extend_immediate_in[14];
			  rotate_immediate_out[21]=extend_immediate_in[13];
			  rotate_immediate_out[20]=extend_immediate_in[12];
			  rotate_immediate_out[19]=extend_immediate_in[11];
			  rotate_immediate_out[18]=extend_immediate_in[10];
			  rotate_immediate_out[17]=extend_immediate_in[9];
			  rotate_immediate_out[16]=extend_immediate_in[8];
			  rotate_immediate_out[15]=extend_immediate_in[7];
			  rotate_immediate_out[14]=extend_immediate_in[6];
			  rotate_immediate_out[13]=extend_immediate_in[5];
			  rotate_immediate_out[12]=extend_immediate_in[4];
			  rotate_immediate_out[11]=extend_immediate_in[3];
			  rotate_immediate_out[10]=extend_immediate_in[2];
			  rotate_immediate_out[9]=extend_immediate_in[1];
			  rotate_immediate_out[8]=extend_immediate_in[0];
			  end
	4'b1101:begin
			  rotate_immediate_out=temp>>26;
			  rotate_immediate_out[31]=extend_immediate_in[25];
			  rotate_immediate_out[30]=extend_immediate_in[24];
			  rotate_immediate_out[29]=extend_immediate_in[23];
			  rotate_immediate_out[28]=extend_immediate_in[22];
			  rotate_immediate_out[27]=extend_immediate_in[21];
			  rotate_immediate_out[26]=extend_immediate_in[20];
			  rotate_immediate_out[25]=extend_immediate_in[19];
			  rotate_immediate_out[24]=extend_immediate_in[18];
			  rotate_immediate_out[23]=extend_immediate_in[17];
			  rotate_immediate_out[22]=extend_immediate_in[16];
			  rotate_immediate_out[21]=extend_immediate_in[15];
			  rotate_immediate_out[20]=extend_immediate_in[14];
			  rotate_immediate_out[19]=extend_immediate_in[13];
			  rotate_immediate_out[18]=extend_immediate_in[12];
			  rotate_immediate_out[17]=extend_immediate_in[11];
			  rotate_immediate_out[16]=extend_immediate_in[10];
			  rotate_immediate_out[15]=extend_immediate_in[9];
			  rotate_immediate_out[14]=extend_immediate_in[8];
			  rotate_immediate_out[13]=extend_immediate_in[7];
			  rotate_immediate_out[12]=extend_immediate_in[6];
			  rotate_immediate_out[11]=extend_immediate_in[5];
			  rotate_immediate_out[10]=extend_immediate_in[4];
			  rotate_immediate_out[9]=extend_immediate_in[3];
			  rotate_immediate_out[8]=extend_immediate_in[2];
			  rotate_immediate_out[7]=extend_immediate_in[1];
			  rotate_immediate_out[6]=extend_immediate_in[0];
			  end
	4'b1110:begin
			  rotate_immediate_out=temp>>28;
			  rotate_immediate_out[31]=extend_immediate_in[27];
			  rotate_immediate_out[30]=extend_immediate_in[26];
			  rotate_immediate_out[29]=extend_immediate_in[25];
			  rotate_immediate_out[28]=extend_immediate_in[24];
			  rotate_immediate_out[27]=extend_immediate_in[23];
			  rotate_immediate_out[26]=extend_immediate_in[22];
			  rotate_immediate_out[25]=extend_immediate_in[21];
			  rotate_immediate_out[24]=extend_immediate_in[20];
			  rotate_immediate_out[23]=extend_immediate_in[19];
			  rotate_immediate_out[22]=extend_immediate_in[18];
			  rotate_immediate_out[21]=extend_immediate_in[17];
			  rotate_immediate_out[20]=extend_immediate_in[16];
			  rotate_immediate_out[19]=extend_immediate_in[15];
			  rotate_immediate_out[18]=extend_immediate_in[14];
			  rotate_immediate_out[17]=extend_immediate_in[13];
			  rotate_immediate_out[16]=extend_immediate_in[12];
			  rotate_immediate_out[15]=extend_immediate_in[11];
			  rotate_immediate_out[14]=extend_immediate_in[10];
			  rotate_immediate_out[13]=extend_immediate_in[9];
			  rotate_immediate_out[12]=extend_immediate_in[8];
			  rotate_immediate_out[11]=extend_immediate_in[7];
			  rotate_immediate_out[10]=extend_immediate_in[6];
			  rotate_immediate_out[9]=extend_immediate_in[5];
			  rotate_immediate_out[8]=extend_immediate_in[4];
			  rotate_immediate_out[7]=extend_immediate_in[3];
			  rotate_immediate_out[6]=extend_immediate_in[2];
			  rotate_immediate_out[5]=extend_immediate_in[1];
			  rotate_immediate_out[4]=extend_immediate_in[0];
			  end
	4'b1111:begin
			  rotate_immediate_out=temp>>30;
			  rotate_immediate_out[31]=extend_immediate_in[29];
			  rotate_immediate_out[30]=extend_immediate_in[28];
			  rotate_immediate_out[29]=extend_immediate_in[27];
			  rotate_immediate_out[28]=extend_immediate_in[26];
			  rotate_immediate_out[27]=extend_immediate_in[25];
			  rotate_immediate_out[26]=extend_immediate_in[24];
			  rotate_immediate_out[25]=extend_immediate_in[23];
			  rotate_immediate_out[24]=extend_immediate_in[22];
			  rotate_immediate_out[23]=extend_immediate_in[21];
			  rotate_immediate_out[22]=extend_immediate_in[20];
			  rotate_immediate_out[21]=extend_immediate_in[19];
			  rotate_immediate_out[20]=extend_immediate_in[18];
			  rotate_immediate_out[19]=extend_immediate_in[17];
			  rotate_immediate_out[18]=extend_immediate_in[16];
			  rotate_immediate_out[17]=extend_immediate_in[15];
			  rotate_immediate_out[16]=extend_immediate_in[14];
			  rotate_immediate_out[15]=extend_immediate_in[13];
			  rotate_immediate_out[14]=extend_immediate_in[12];
			  rotate_immediate_out[13]=extend_immediate_in[11];
			  rotate_immediate_out[12]=extend_immediate_in[10];
			  rotate_immediate_out[11]=extend_immediate_in[9];
			  rotate_immediate_out[10]=extend_immediate_in[8];
			  rotate_immediate_out[9]=extend_immediate_in[7];
			  rotate_immediate_out[8]=extend_immediate_in[6];
			  rotate_immediate_out[7]=extend_immediate_in[5];
			  rotate_immediate_out[6]=extend_immediate_in[4];
			  rotate_immediate_out[5]=extend_immediate_in[3];
			  rotate_immediate_out[4]=extend_immediate_in[2];
			  rotate_immediate_out[3]=extend_immediate_in[1];
			  rotate_immediate_out[2]=extend_immediate_in[0];
			  end
	endcase

end

endmodule